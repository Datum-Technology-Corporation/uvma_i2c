// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_I2C_ST_TDEFS_SV__
`define __UVMT_I2C_ST_TDEFS_SV__





`endif // __UVMT_I2C_ST_TDEFS_SV__