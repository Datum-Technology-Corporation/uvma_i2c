// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_I2C_ST_MACROS_SV__
`define __UVMT_I2C_ST_MACROS_SV__





`endif // __UVMT_I2C_ST_MACROS_SV__