// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_I2C_ST_CONSTANTS_SV__
`define __UVME_I2C_ST_CONSTANTS_SV__


const int unsigned uvme_i2c_st_rand_stim_default_num_seq_items =    10; ///< Default number of Sequence Items generated by uvme_i2c_st_rand_stim_vseq_c in each direction.
const int unsigned uvme_i2c_st_rand_stim_sqr_priority          = 1_000; ///< Sequencer priority for uvme_i2c_st_rand_stim_vseq_c Sequence Items.


`endif // __UVME_I2C_ST_CONSTANTS_SV__