// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_I2C_ST_MACROS_SV__
`define __UVME_I2C_ST_MACROS_SV__


// Add preprocessor macros here
// Ex: `ifndef UVME_${name_uppercase}_ST_ABC
//        `define UVME_${name_uppercase}_ST_ABC 32
//     `endif


`endif // __UVME_I2C_ST_MACROS_SV__