// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_I2C_MACROS_SV__
`define __UVMA_I2C_MACROS_SV__


`define UVMA_I2C_C2T_DRV_SEQ_ITEM_PRI  100
`define UVMA_I2C_T2C_DRV_SEQ_ITEM_PRI  100
`define UVMA_I2C_IDLE_SEQ_ITEM_PRI  1


`endif // __UVMA_I2C_MACROS_SV__